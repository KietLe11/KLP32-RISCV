module RV32I(clk);

input wire clk;

endmodule