`timescale 1 ns/1 ps
module register32_tb();

    parameter n = 32;
    reg [n-1:0] write_data

endmodule