module KLP32V1(clk);

input wire clk;

endmodule